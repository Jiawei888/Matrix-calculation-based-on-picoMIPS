//----------------------------------------------------- 
// File Name : alucodes.sv
// FuncRon
// Author: tjk
// Last rev. 23 Oct 12 //----------------------------------------------------- //
`define RADD 3'b010
`define RSUB 3'b011
`define MUL 3'b111