//----------------------------------------------------- 
// File Name : opcodes.sv
// FuncRon
// Author: ljw
// Last rev. 16 Febr 20 //----------------------------------------------------- //
`define NOP 6'b000000
`define ADD 6'b000010
`define SUB 6'b000011
`define ADDI 6'b001010
`define SUBI 6'b001011
`define MUL 6'b010111

